module top(
in
)