module top();
    
endmodule //top
