module mux