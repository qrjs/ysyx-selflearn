module top(
    input []
);
    
endmodule //top

