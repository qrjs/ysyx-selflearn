module mux41(
    input [1:0] sel,
    
)