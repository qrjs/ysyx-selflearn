module top(
    input [7:0]
);
    
endmodule //top

