module top(
    input [7:0]x,
    input en,
    i
);
    
endmodule //top

