module moduleName();
    
endmodule //moduleName
