module top(
    input [3:0] A,B,
    IN
);
    
endmodule //top
