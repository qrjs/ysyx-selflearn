module top(
    
)