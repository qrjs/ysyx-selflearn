module mux41(
    input [1:0] sel,
    input [1]
)