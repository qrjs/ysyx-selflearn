module top(
    input [3:0] a,
    input [2:0] alu_ch
    output [3:0] f
);
    
endmodule //top
