module top(
    
);
    
endmodule //top

