module mux21(
    input
)