module top(
    input [3:0] A,B,
    input [2:0] alu_ch
    output [3:0] $fclose();
);
    
endmodule //top
