module top(
    input [7]
)