module moduleName (
    input      clk,
    input      rst,
    
);
    
endmodule //moduleName
