module top(
    input [7:0] din,
    input [2:0] shamt,
    input LR,
    input AL,
    output reg [7:0] dout
);
wire w0,w1,w2,w3,w4,w5,w6,w7,w8,w9,w10,w11,w12,w13,w14,w15,w16;

// 修改实例名称
mux21 u_0_1(.sel(AL), .x0(0), .x1(din[7]), .f(w0));
mux41 u_1_1(.sel({LR, shamt[0]}), .x0(din[7]), .x1(w0), .x2(din[7]), .x3(din[6]), .f(w1));
mux41 u_2_1(.sel({LR, shamt[0]}), .x0(din[6]), .x1(din[7]), .x2(din[6]), .x3(din[5]), .f(w2));
mux41 u_3_1(.sel({LR, shamt[0]}), .x0(din[5]), .x1(din[6]), .x2(din[5]), .x3(din[4]), .f(w3));
mux41 u_4_1(.sel({LR, shamt[0]}), .x0(din[4]), .x1(din[5]), .x2(din[4]), .x3(din[3]), .f(w4));
mux41 u_5_1(.sel({LR, shamt[0]}), .x0(din[3]), .x1(din[4]), .x2(din[3]), .x3(din[2]), .f(w5));
mux41 u_6_1(.sel({LR, shamt[0]}), .x0(din[2]), .x1(din[3]), .x2(din[2]), .x3(din[1]), .f(w6));
mux41 u_7_1(.sel({LR, shamt[0]}), .x0(din[1]), .x1(din[2]), .x2(din[1]), .x3(din[0]), .f(w7));
mux41 u_8_1(.sel({LR, shamt[0]}), .x0(din[0]), .x1(din[1]), .x2(din[0]), .x3(0), .f(w8));

mux41 u_1_2(.sel({LR, shamt[1]}), .x0(w1), .x1(w0), .x2(w1), .x3(w3), .f(w9));
mux41 u_2_2(.sel({LR, shamt[1]}), .x0(w2), .x1(w0), .x2(w2), .x3(w4), .f(w10));
mux41 u_3_2(.sel({LR, shamt[1]}), .x0(w3), .x1(w1), .x2(w3), .x3(w5), .f(w11));
mux41 u_4_2(.sel({LR, shamt[1]}), .x0(w4), .x1(w2), .x2(w4), .x3(w6), .f(w12));
mux41 u_5_2(.sel({LR, shamt[1]}), .x0(w5), .x1(w3), .x2(w5), .x3(w7), .f(w13));
mux41 u_6_2(.sel({LR, shamt[1]}), .x0(w6), .x1(w4), .x2(w6), .x3(w8), .f(w14));
mux41 u_7_2(.sel({LR, shamt[1]}), .x0(w7), .x1(w5), .x2(w7), .x3(0), .f(w15));
mux41 u_8_2(.sel({LR, shamt[1]}), .x0(w8), .x1(w6), .x2(w8), .x3(0), .f(w16));

mux41 u_1_3(.sel({LR, shamt[2]}), .x0(w9), .x1(w0), .x2(w9), .x3(w13), .f(dout[7]));
mux41 u_2_3(.sel({LR, shamt[2]}), .x0(w10), .x1(w0), .x2(w10), .x3(w14), .f(dout[6]));
mux41 u_3_3(.sel({LR, shamt[2]}), .x0(w11), .x1(w0), .x2(w11), .x3(w15), .f(dout[5]));
mux41 u_4_3(.sel({LR, shamt[2]}), .x0(w12), .x1(w0), .x2(w12), .x3(w16), .f(dout[4]));
mux41 u_5_3(.sel({LR, shamt[2]}), .x0(w13), .x1(w9), .x2(w13), .x3(0), .f(dout[3]));
mux41 u_6_3(.sel({LR, shamt[2]}), .x0(w14), .x1(w10), .x2(w14), .x3(0), .f(dout[2]));
mux41 u_7_3(.sel({LR, shamt[2]}), .x0(w15), .x1(w11), .x2(w15), .x3(0), .f(dout[1]));
mux41 u_8_3(.sel({LR, shamt[2]}), .x0(w16), .x1(w12), .x2(w16), .x3(0), .f(dout[0]));

endmodule
