module top(
    input [7:0]x,
    input en,
    output reg vx,
    output reg [2:0] y,
    output reg 
);
    
endmodule //top

