module top(
    input [7:0] din,
    input []
)