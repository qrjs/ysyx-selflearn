module mux21(
    input sel
)