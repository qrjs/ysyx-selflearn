module top(
    input [7:0] din,
    input [2:0 ]
)