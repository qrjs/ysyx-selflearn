module top(
    input [3:0] A,B,
    in
);
    
endmodule //top
