module top(
    input [7:0]x,
    input en,
    output 
);
    
endmodule //top

