module mux41(

)