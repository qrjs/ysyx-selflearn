module top(
    input [3:0] A,B,
    input []
);
    
endmodule //top
