module top(
    input [7:0]x,
    
);
    
endmodule //top

