module top(
    
);
    
endmodule //top
