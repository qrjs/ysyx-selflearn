module top(
    input [7:0]x,
    input en,
    output reg vx,
    output reg 
);
    
endmodule //top

