module top(
    input [7:0] din,
    input [2:0] shamt,
    input LR,
    input 
)