module mux41(
    input [1:0] sel,
    input [1:0] x0,x2,x3,x4,
    output reg [1:0] f
);
always@(*)begin
    case(sel)
    
end
