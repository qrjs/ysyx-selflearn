module mux21(
    input sel,
    input x0,x1,
    output reg f
);
always