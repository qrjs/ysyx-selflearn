module top(
    input [3:0] a,b,
    input [2:0] alu_ch
    output [3:0] alu_f,
    output zero_f,over_f,cin_f
);
    
endmodule //top
